Testing for initial commit github
